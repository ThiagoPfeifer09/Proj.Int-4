module cache_dados (
    input logic clk,
    input logic reset,  // antes era rst

    input logic [31:0] address,
    input logic [63:0] write_data,
    input logic mem_read,
    input logic mem_write,

    output logic [63:0] read_data,  // antes era data_out
    output logic miss,              // antes era ready

    // interface com a memória principal
    output logic [31:0] mem_address,
    output logic [63:0] mem_write_data,
    input logic [127:0] mem_block_read_data,
    input logic mem_ready,
    output logic mem_read_out,
    output logic mem_write_out
);

    typedef enum logic [1:0] {
        IDLE,
        MISS
    } state_t;

    state_t state;

    typedef struct packed {
        logic valid;
        logic [24:0] tag;
        logic [127:0] data;
    } cache_line_t;

    cache_line_t cache [0:3];

    logic [1:0] index;
    logic [24:0] tag;
    logic [3:0] offset;

    assign index = address[3:2];
    assign tag = address[31:7];
    assign offset = address[6:3];

    always_ff @(posedge clk or posedge reset) begin
        if (reset) begin
            state <= IDLE;
            miss <= 0;
            read_data <= 0;
            mem_read_out <= 0;
            mem_write_out <= 0;
            for (int i = 0; i < 4; i++) begin
                cache[i].valid <= 0;
                cache[i].tag <= 0;
                cache[i].data <= 0;
            end
        end else begin
            case (state)
                IDLE: begin
                    mem_read_out <= 0;
                    mem_write_out <= 0;
                    miss <= 0;

                    if (mem_read && !mem_write) begin
                        if (cache[index].valid && cache[index].tag == tag) begin
                            // HIT leitura
                            case (offset[3:3])
                                1'b0: read_data <= cache[index].data[63:0];
                                1'b1: read_data <= cache[index].data[127:64];
                            endcase
                            miss <= 1;
                        end else begin
                            // MISS leitura
                            mem_address <= {address[31:4], 4'b0000};
                            mem_read_out <= 1;
                            state <= MISS;
                        end
                    end else if (mem_write) begin
                        // Escrita direta (write-through)
                        mem_address <= address;
                        mem_write_data <= write_data;
                        mem_write_out <= 1;

                        // Atualiza cache se HIT
                        if (cache[index].valid && cache[index].tag == tag) begin
                            if (offset[3:3] == 1'b0) begin
                                cache[index].data[63:0] <= write_data;
                                read_data <= write_data;
                            end else begin
                                cache[index].data[127:64] <= write_data;
                                read_data <= write_data;
                            end
                        end

                        miss <= 1;
                    end
                end

                MISS: begin
                    if (mem_ready) begin
                        // Refill da cache
                        cache[index].valid <= 1;
                        cache[index].tag <= tag;
                        cache[index].data <= mem_block_read_data;

                        // Entrega o dado ao processador
                        case (offset[3:3])
                            1'b0: read_data <= mem_block_read_data[63:0];
                            1'b1: read_data <= mem_block_read_data[127:64];
                        endcase

                        miss <= 1;
                        state <= IDLE;
                    end
                end
            endcase
        end
    end
endmodule
