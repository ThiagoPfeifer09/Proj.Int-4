module riscv_pipeline (input wire clk, input wire rst);
    wire [31:0] if_id_pc_out, if_id_pc_4_out, if_id_instr_out;
    wire [31:0] id_ex_pc_out, id_ex_pc_4_out, id_ex_rs1_data_out, id_ex_rs2_data_out, id_ex_imm_out;
    wire [4:0]  id_ex_rd_out, id_ex_rs1_out, id_ex_rs2_out;
    wire [2:0]  id_ex_funct3_out; wire [6:0]  id_ex_funct7_out, id_ex_opcode_out;
    wire [31:0] ex_mem_pc, ex_mem_pc_4, ex_mem_alu_result, ex_mem_rs2_data;
    wire [4:0]  ex_mem_rd; wire [2:0]  ex_mem_funct3; wire [6:0]  ex_mem_opcode;
    wire        ex_mem_mem_write_en, ex_mem_mem_read_en, ex_mem_reg_write_en;
    wire [1:0]  ex_mem_mem_to_reg_sel;
    wire [31:0] mem_wb_pc_4, mem_wb_alu_result, mem_wb_mem_read_data;
    wire [4:0]  mem_wb_rd; wire        mem_wb_reg_write_en; wire [1:0]  mem_wb_mem_to_reg_sel;
    wire [31:0] wb_to_rf_reg_write_data;
    wire        pc_write_en, if_id_write_en;
    wire [31:0] branch_target_from_ex; wire        branch_taken_from_ex;
    wire [31:0] mem_addr_to_dm, mem_write_data_to_dm, mem_read_data_from_dm;
    wire        mem_write_byte_en_to_dm, mem_write_half_en_to_dm, mem_write_word_en_to_dm;

    if_stage u_if_stage ( .clk(clk), .rst(rst), .branch_target_in(branch_target_from_ex), .branch_taken_in(branch_taken_from_ex), .pc_write_en_in(pc_write_en), .if_id_write_en_in(if_id_write_en), .if_id_pc_out(if_id_pc_out), .if_id_pc_4_out(if_id_pc_4_out), .if_id_instr_out(if_id_instr_out) );
    id_stage u_id_stage ( .clk(clk), .rst(rst), .if_id_pc_in(if_id_pc_out), .if_id_pc_4_in(if_id_pc_4_out), .if_id_instr_in(if_id_instr_out), .ex_mem_mem_read_en_in(ex_mem_mem_read_en), .ex_mem_rd_in(ex_mem_rd), .branch_taken_from_ex_in(branch_taken_from_ex), .mem_wb_reg_write_en_in(mem_wb_reg_write_en), .mem_wb_rd_in(mem_wb_rd), .mem_wb_write_data_in(wb_to_rf_reg_write_data), .pc_write_en_out(pc_write_en), .if_id_write_en_out(if_id_write_en), .id_ex_pc_out(id_ex_pc_out), .id_ex_pc_4_out(id_ex_pc_4_out), .id_ex_rs1_data_out(id_ex_rs1_data_out), .id_ex_rs2_data_out(id_ex_rs2_data_out), .id_ex_rd_out(id_ex_rd_out), .id_ex_rs1_out(id_ex_rs1_out), .id_ex_rs2_out(id_ex_rs2_out), .id_ex_funct3_out(id_ex_funct3_out), .id_ex_funct7_out(id_ex_funct7_out), .id_ex_opcode_out(id_ex_opcode_out), .id_ex_imm_out(id_ex_imm_out) );
    ex_stage u_ex_stage ( .clk(clk), .rst(rst), .id_ex_pc(id_ex_pc_out), .id_ex_pc_4(id_ex_pc_4_out), .id_ex_rs1_data(id_ex_rs1_data_out), .id_ex_rs2_data(id_ex_rs2_data_out), .id_ex_rd(id_ex_rd_out), .id_ex_rs1(id_ex_rs1_out), .id_ex_rs2(id_ex_rs2_out), .id_ex_funct3(id_ex_funct3_out), .id_ex_funct7(id_ex_funct7_out), .id_ex_opcode(id_ex_opcode_out), .id_ex_imm(id_ex_imm_out), .ex_mem_rd_in(ex_mem_rd), .ex_mem_reg_write_en_in(ex_mem_reg_write_en), .ex_mem_alu_result_in(ex_mem_alu_result), .mem_wb_rd_in(mem_wb_rd), .mem_wb_reg_write_en_in(mem_wb_reg_write_en), .mem_wb_write_data_in(wb_to_rf_reg_write_data), .ex_mem_pc(ex_mem_pc), .ex_mem_pc_4(ex_mem_pc_4), .ex_mem_alu_result(ex_mem_alu_result), .ex_mem_rs2_data(ex_mem_rs2_data), .ex_mem_rd(ex_mem_rd), .ex_mem_funct3(ex_mem_funct3), .ex_mem_opcode(ex_mem_opcode), .ex_mem_mem_write_en(ex_mem_mem_write_en), .ex_mem_mem_read_en(ex_mem_mem_read_en), .ex_mem_reg_write_en(ex_mem_reg_write_en), .ex_mem_mem_to_reg_sel(ex_mem_mem_to_reg_sel), .branch_target(branch_target_from_ex), .branch_taken(branch_taken_from_ex) );
    mem_stage u_mem_stage ( .clk(clk), .rst(rst), .ex_mem_pc(ex_mem_pc), .ex_mem_pc_4(ex_mem_pc_4), .ex_mem_alu_result(ex_mem_alu_result), .ex_mem_rs2_data(ex_mem_rs2_data), .ex_mem_rd(ex_mem_rd), .ex_mem_funct3(ex_mem_funct3), .ex_mem_opcode(ex_mem_opcode), .ex_mem_mem_write_en(ex_mem_mem_write_en), .ex_mem_mem_read_en(ex_mem_mem_read_en), .ex_mem_reg_write_en(ex_mem_reg_write_en), .ex_mem_mem_to_reg_sel(ex_mem_mem_to_reg_sel), .mem_addr(mem_addr_to_dm), .mem_write_data(mem_write_data_to_dm), .mem_write_byte_en(mem_write_byte_en_to_dm), .mem_write_half_en(mem_write_half_en_to_dm), .mem_write_word_en(mem_write_word_en_to_dm), .mem_read_data(mem_read_data_from_dm), .mem_wb_pc_4(mem_wb_pc_4), .mem_wb_alu_result(mem_wb_alu_result), .mem_wb_mem_read_data(mem_wb_mem_read_data), .mem_wb_rd(mem_wb_rd), .mem_wb_reg_write_en(mem_wb_reg_write_en), .mem_wb_mem_to_reg_sel(mem_wb_mem_to_reg_sel) );
    wb_stage u_wb_stage ( .clk(clk), .rst(rst), .mem_wb_pc_4(mem_wb_pc_4), .mem_wb_alu_result(mem_wb_alu_result), .mem_wb_mem_read_data(mem_wb_mem_read_data), .mem_wb_rd(mem_wb_rd), .mem_wb_reg_write_en(mem_wb_reg_write_en), .mem_wb_mem_to_reg_sel(mem_wb_mem_to_reg_sel), .reg_write_en_out(), .reg_write_addr_out(), .reg_write_data_out(wb_to_rf_reg_write_data) );
    data_mem u_data_mem ( .clk(clk), .addr(mem_addr_to_dm), .write_data(mem_write_data_to_dm), .read_en(ex_mem_mem_read_en), .write_byte_en(mem_write_byte_en_to_dm), .write_half_en(mem_write_half_en_to_dm), .write_word_en(mem_write_word_en_to_dm), .read_data(mem_read_data_from_dm) );
endmodule